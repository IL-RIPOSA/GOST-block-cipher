library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity s_box_arr is
	port(
	data: in std_logic_vector(31 downto 0);
	data_out: out std_logic_vector(31 downto 0)
	);
end s_box_arr;

architecture s_box_arr_arch of s_box_arr is

type array2D is array (7 downto 0, 0 to 15) of std_logic_vector(3 downto 0);
signal s_array: array2D:=(
		( "0100", "1010", "1001", "0010", "1101", "1000", "0000", "1110", "0110", "1011", "0001", "1100", "0111", "1111", "0101", "0011" ),--MSB
    		( "1110", "1011", "0100", "1100", "0110", "1101", "1111", "1010", "0010", "0011", "1000", "0001", "0000", "0111", "0101", "1001" ),
    		( "0101", "1000", "0001", "1101", "1010", "0011", "0100", "0010", "1110", "1111", "1100", "0111", "0110", "0000", "1001", "1011" ),
    		( "0111", "1101", "1010", "0001", "0000", "1000", "1001", "1111", "1110", "0100", "0110", "1100", "1101", "0010", "0101", "0011" ),
    		( "0110", "1100", "0111", "0001", "0101", "1111", "1101", "1000", "0100", "1010", "1001", "1110", "0000", "0011", "1011", "0010" ),
   		( "0100", "1011", "1010", "0000", "0111", "0010", "0001", "1101", "0011", "0110", "1000", "0101", "1001", "1100", "1111", "1110" ),
   		( "1101", "1011", "0100", "0001", "0011", "1111", "0101", "1001", "0000", "1010", "1110", "0110", "1100", "1000", "0010", "1100" ),
  		( "0001", "1111", "1101", "0000", "0101", "0111", "1010", "0100", "1001", "0010", "0011", "1110", "0110", "1011", "1000", "1100" ) --LSB
		 );

begin
	G1:for i in 0 to 7 generate
		data_out(4*i+3 downto 4*i)<= s_array(i,to_integer(unsigned(data(4*i+3 downto 4*i))));
	end generate;

end s_box_arr_arch;